module top (output [7:0] LED);

	assign LED= 8'b11111111;

endmodule
